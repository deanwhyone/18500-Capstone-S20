/*
 * 18500 Capstone S20
 * Eric Chen, Alton Olsen, Deanyone Su
 *
 */
 `default_nettype none

module Sender
	import NetworkPkg::*,
		   DisplayPkg::*;
(

);

endmodule // Sender