/*
 * 18500 Capstone S20
 * Eric Chen, Alton Olsen, Deanyone Su
 * Serial data sender for single data wire
 */
 `default_nettype none

module DataSender
	import NetworkPkg::*,
		   DisplayPkg::*;
(

);

endmodule // DataSender