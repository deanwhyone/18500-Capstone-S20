/*
 * 18500 Capstone S20
 * Eric Chen, Alton Olsen, Deanyone Su
 * Serial data sender for handshake wire
 */
 `default_nettype none

module HandshakeSender
	import NetworkPkg::*,
		   DisplayPkg::*;
(

);

endmodule // HandshakeSender